//Subject:     LAB4
//--------------------------------------------------------------------------------
//Version:     1
//--------------------------------------------------------------------------------
//Writer:      高鈺鴻
//----------------------------------------------
//Date: 2022/5/25
//----------------------------------------------
//Description:
//--------------------------------------------------------------------------------

module Shift_Left_Two_32(
    data_i,
    data_o
  );

  //I/O ports
  input [32-1:0] data_i;
  output [32-1:0] data_o;

  //shift left 2
  assign data_o = {data_i[30-1:0],2'b00};
endmodule
