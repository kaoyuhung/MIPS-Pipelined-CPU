//Subject:     LAB4
//--------------------------------------------------------------------------------
//Version:     1
//--------------------------------------------------------------------------------
//Writer:      高鈺鴻
//----------------------------------------------
//Date: 2022/5/25
//----------------------------------------------
//Description:
//--------------------------------------------------------------------------------

module Sign_Extend(
    data_i,
    data_o
  );

  //I/O ports
  input   [16-1:0] data_i;
  output  [32-1:0] data_o;

  //Internal Signals
  reg     [32-1:0] data_o;

  //Sign extended
  always @(*)
  begin
    data_o <= {{16{data_i[16-1]}},data_i};
  end
endmodule

